module power

// Simple tests for the power function
fn test_power() {
	assert power(2.0, 3.0) == 8.0
	assert power(5.0, 3.0) == 125.0
}
